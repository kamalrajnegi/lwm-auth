/*

Designed By:
Kamal Raj (kamal@kamalraj.in)
*/
module demo_puf(
    clk,
    challenge,
    response,
);


//puf code will be added in the future


endmodule