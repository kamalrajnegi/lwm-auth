/*
Designed By:
Kamal Raj (kamal@kamalraj.in)
*/
module lwm_auth_top(
    clk,
    enable,
    tx,
    tx,
    done
);


//the design will be added here in the future


endmodule