/*
Designed By:
Kamal Raj (kamal@kamalraj.in)
*/
module ascon(
    clk,
    start,
    key,
    data_in,
    data_out,
    address_in,
    address_out
);


// ASCON design will be added here in the future


endmodule